`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:25:34 11/17/2022 
// Design Name: 
// Module Name:    controllBuzz 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module controllBuzz(switch,notes);
	input [6:0] switch
	input [6:0] notes
	output speaker
	reg [6:0] currentSW
	
	always @(posedge clk) begin
		
			
	
endmodule
